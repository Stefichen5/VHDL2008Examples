package packGenerateType is
	type aThingToGenerate is (ComponentA, ComponentB, ComponentC, ComponentD);
end package packGenerateType;

package body packGenerateType is
	
end package body packGenerateType;
